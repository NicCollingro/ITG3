module top_level();
    reg clk = 1;
    always #1 = ~clk;
    reg g,y,r;
    reg [2,0] cnt;
    




endmodule