// TOPLEVEL oberstes Modul
module test1 ;


endmodule;


// TESTBENCH