module top_level(CLOCK_50,GPIO_023,GPIO_021,
 GPIO_019,GPIO_017, GPIO_015,GPIO_013,GPIO_011);
input CLOCK_50, ;

always

endmodule

module keypad(input clk; output reg [3:0] keycode,
input [2:0] cols, output reg [3:0] rows);


endmodule