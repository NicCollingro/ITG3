module I2C_master (input wire sda, output wire scl, input wire send, output wire busy,
input wire [6:0] addr, input wire [7:0] data , input wire rw);



endmodule