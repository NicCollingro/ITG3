../../src_common/symbols.vh