`define BASECLK CLOCK_HALF // Pixel Clock
`define HRES 640 // horizontal resolution
`define HSRT 656 // hsync pulse start
`define HEND 752 // hsync pulse end
`define HTOT 800 // line end
`define VRES 480 // vertical resolution
`define VSRT 490 // vsync pulse start
`define VEND 492 // vsync pulse end
`define VTOT 525 // frame end