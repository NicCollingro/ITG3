module control(input wire[7:0] state, input wire [2:0] operand1, 
input wire [2:0]operand2, input wire flag_carry, input wire flag_zero,
output wire c_ii, c_ci, c_co, c_cs, c_rfi, c_rfo, c_eo, c_ee, c_mi, 
c_ro, c_ri, c_so, c_sd, c_si, c_halt);



endmodule