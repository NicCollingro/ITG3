module computer (CLOCK_50);
inout wire data_bus

endmodule