module top_level();
    reg clk = 1;
    always #1 = ~clk;
    reg g,y,r;
    




endmodule